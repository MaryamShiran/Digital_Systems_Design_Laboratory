library verilog;
use verilog.vl_types.all;
entity TB_FI is
end TB_FI;
