library verilog;
use verilog.vl_types.all;
entity TB_Booth is
end TB_Booth;
